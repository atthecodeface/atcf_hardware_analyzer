/** @copyright (C) 2020,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   analyzer_target.cdl
 * @brief  Standard target for the analyzer bus
 *

 */

/*a Includes
 */
include "analyzer.h"
include "analyzer_modules.h"

/*a Module
 */
/*m analyzer_target_stub
 *
 * Stub for the logic analyzer bus with no source (to plug muxes)
 *
 */
module analyzer_target_stub( clock clk,
                        input bit reset_n,

                        input  t_analyzer_mst  analyzer_mst,
                        output t_analyzer_tgt  analyzer_tgt
    )
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;

    /*b APB interface state  */
    net t_analyzer_tgt analyzer_tgt;
    clocked t_analyzer_data4 analyzer_data = {*=0};

    /*b Blah */
    blah : {
        analyzer_data <= {*=0};
        analyzer_target stub( clk<-clk, reset_n<=reset_n,
                              analyzer_mst <= analyzer_mst,
                              analyzer_tgt => analyzer_tgt,
                              // analyzer_ctl =>
                              analyzer_data <= analyzer_data );
    }

    /*b All done */
}
