/*a Includes
 */
include "apb::apb.h"
include "analyzer.h"
include "std::tech_sync.h"
include "std::srams.h"

/*a Constants
 */
constant integer analyzer_signal_width = 32;
constant integer analyzer_trigger_signal_width = 32;
constant integer analyzer_trigger_counter_width = 16;
constant integer analyzer_trigger_depth_log = 2;
constant integer analyzer_trigger_depth = 4;
constant integer analyzer_ram_depth_log = 11; // 2048 by 32 for the RAM sounds good

/*a Types */
/*t t_analyzer_action
 */
typedef enum [3]
{
    analyzer_action_idle,                           // H Store nothing, and do not touch counter
    analyzer_action_reset_counter,                  // L Store nothing, and reset counter to 1, stay in current stage
    analyzer_action_store_signal_and_transition,    // M Store signal value and transition immediately
    analyzer_action_store_signal_and_reside,        // H Store signal value and transition if counter matches residence time
    analyzer_action_store_time_and_reside,          // L Store time of occurrence (cycles since trigger_reset went away) and trigger signals, transition if counter matches residence time
    analyzer_action_store_time_and_transition,      // H Store time of occurrence (cycles since trigger_reset went away) and trigger signals and transition
    analyzer_action_store_residence_and_transition, // M Store residence time and transition
    analyzer_action_end,                            // H Store nothing, disable trace
//    analyzer_action_compress,
} t_analyzer_action;

/*t t_trigger_store_type
 */
typedef enum [2]
{
    trigger_store_type_none,
    trigger_store_type_signal,
    trigger_store_type_time,
    trigger_store_type_residence
} t_trigger_store_type;

/*t t_analyzer_trigger
 */
typedef struct
{
    bit[analyzer_trigger_signal_width] mask     "Mask for incoming signal bits";
    bit[analyzer_trigger_signal_width] compare  "Value the masked signal should be to match";
    bit[analyzer_trigger_counter_width] counter "Number of cycles that the masked signal should match; ==0 means only leave if false";
    bit[analyzer_trigger_depth_log] if_false    "State to enter if masked value does not match";
    bit[analyzer_trigger_depth_log] if_true     "State to enter if masked value matched for cycle given by 'counter'";
    t_analyzer_action action_if_true "Action to take whilst in this state and true";
    t_analyzer_action action_if_false "Action to take whilst in this state and true";
} t_analyzer_trigger;

/*t t_apb_address
 * APB address map, used to decode paddr
 */
typedef enum [4] {
    apb_address_config      = 0,
    apb_address_trigger     = 1,
    apb_address_mask        = 2,
    apb_address_compare     = 3,
    apb_address_mux_control = 4,
    apb_address_trace_data  = 8,
} t_apb_address;

/*t t_access
 * APB access that is in progress; a decode of psel and paddr
 */
typedef enum [3] {
    access_none                     "No access being performed",
    access_write_config             "Writing config",
    access_write_trigger            "Write trigger transition and counter",
    access_write_mask               "Write trigger mask",
    access_write_compare            "Write trigger compare",
    access_write_mux_control        "Write analyzer mux control",
    access_read_status              "Read status",
    access_read_trace_data          "Read trace data",
} t_access;

/*t t_apb_combs */
typedef struct {
    bit unused;
} t_apb_combs;

/*t t_analyzer_control_fsm */
typedef fsm {
    actl_idle;
    actl_enable;
    actl_data;
} t_analyzer_control_fsm;

/*t t_analyzer_control */
typedef struct {
    bit enable;
    bit write_data;
    bit[3]  nybbles;
    bit[24] data;
    t_analyzer_control_fsm state;
} t_analyzer_control;

/*t t_apb_state */
typedef struct {
    t_analyzer_control control;
    t_access access;
    bit last_valid_sync;
    bit trace_req;
} t_apb_state;

/*a Module
 */
module apb_target_simple_analyzer( clock clk,

                                   input bit reset_n,

                                   input  t_apb_request  apb_request  "APB request",
                                   output t_apb_response apb_response "APB response",

                                   input t_timer_value timer_value,
                                   input t_analyzer_data4 analyzer_data
    )
"""
"""

{
    /*b Default clock and reset
     */
    default clock analyzer_clock;
    default reset active_low reset_n;

    /*b Outputs for the async trace read interface
     */
    clocked clock async_trace_read_clock bit async_trace_valid_out = 0;
    clocked clock async_trace_read_clock bit[analyzer_signal_width] async_trace_out = 0;

    /*b APB interface
     */
    clocked clock apb_clock bit apb_trigger_reset = 0;
    clocked clock apb_clock bit apb_trigger_enable = 0;
    clocked clock apb_clock bit[analyzer_trigger_depth_log] apb_trigger_stage = 0;
    clocked clock apb_clock bit apb_trace_readback = 0; // asserted if APB should read data from circular buffer
    clocked clock apb_clock bit[32] apb_trace_data = 0;
    clocked clock apb_clock bit apb_trace_valid = 0;
    comb bit apb_read_trace;

    /*b Synchronize and read out of FIFO to APB
     */
    net bit apb_valid_sync;
    //comb    t_apb_combs  apb_combs;
    clocked clock apb_clock t_apb_state apb_state = {*=0};

    /*b Trigger
     */
    clocked clock apb_clock t_analyzer_trigger[analyzer_trigger_depth] trigger = { { mask=0, compare=0, counter=0, if_false=0, if_true=0, action_if_false=analyzer_action_idle, action_if_true=analyzer_action_idle } };
    clocked bit trigger_reset = 0;
    clocked bit trigger_enable = 0;
    clocked bit trigger_done = 0;
    clocked bit trigger_circular = 0;
    clocked bit[analyzer_trigger_depth_log] trigger_stage = 0;
    clocked bit[analyzer_trigger_counter_width] trigger_residence = 1;
    clocked bit[24] trigger_time=0;
    comb bit[analyzer_trigger_signal_width] trigger_mask;
    comb bit[analyzer_trigger_signal_width] trigger_compare;
    comb bit trigger_match;
    comb t_analyzer_action trigger_action;
    comb bit trigger_transition;
    comb bit trigger_hold_counter;
    comb bit trigger_reset_counter;
    comb bit trigger_residence_expired;
    comb bit action_trigger_end;
    comb t_trigger_store_type trigger_store_type;

    /*b Register incoming data and store in FIFO
     */
    clocked t_analyzer_tgt analyzer_tgt_r =  {*=0};
    clocked t_analyzer_mst analyzer_mst = {*=0};
    comb bit[analyzer_signal_width] buffered_input;
    clocked bit[analyzer_ram_depth_log] write_ptr = 0;

    /*b Read out of FIFO
     */
    clocked bit[analyzer_ram_depth_log] read_ptr = 0;
    clocked bit fifo_reading = 0;
    net bit[analyzer_signal_width] fifo_read_data;
    clocked bit[analyzer_signal_width] buffered_read_data=0;
    comb bit fifo_empty;
    comb bit fifo_full;
    comb bit fifo_write;
    comb bit[analyzer_signal_width] fifo_write_data;
    comb bit fifo_read;
    comb bit fifo_end_trigger;
    comb bit fifo_inc_read_ptr;
    clocked bit int_req_sync_0 = 0;
    clocked bit int_req_sync_1 = 0;
    clocked bit valid = 0;

    /*b Synchronize and read out of FIFO to our async read port
     */
    net bit async_out_valid_sync;
    clocked clock async_trace_read_clock bit async_out_last_valid_sync = 0;
    clocked clock async_trace_read_clock bit async_trace_req = 0;

    /*b Trigger and trace ram
     */
    trigger_and_trace_ram "Trigger and trace RAM": {
        

        analyzer_trigger_simple trigger( clk <- clk,
                                         reset_n <= reset_n,
                                         din <= analyzer_data,
                                         dout => trigger_dout,
                                         trace_op => trace_op,
                                         timer_value <= timer_value,
                                         trigger_cfg <= trigger_cfg
            );
        analyzer_trace_ram trace( clk <- clk,
                                  reset_n <= reset_n,

                                  trace_op <= trace_op,
                                  din <= trigger_dout,
                                  fifo_status_l => trace_fifo_status[0],
                                  fifo_status_h => trace_fifo_status[1],

                                  trace_req <= trace_req,
                                  trace_resp => trace_resp,
                                  trace_cfg <= trace_cfg
            );
        )
        analyzer_tgt_r <= analyzer_tgt;
        buffered_input = analyzer_tgt_r.data.data[32;0]; // for now...
        full_switch (apb_state.control.state) {
        case actl_idle: {
            analyzer_mst.select <= 0;
            if (apb_state.control.enable  && !analyzer_mst.enable) {
                apb_state.control.state <= actl_enable;
            }
            if (!apb_state.control.enable && analyzer_mst.enable) {
                analyzer_mst <= {*=0};
            }
            if (apb_state.control.write_data) {
                apb_state.control.state <= actl_data;
            }
        }
        case actl_enable: {
            analyzer_mst.enable <= 1;
            if (apb_state.control.data==0) {
                analyzer_mst.select <= 1;
                apb_state.control.state <= actl_idle;
            } else {
                apb_state.control.data <= apb_state.control.data - 1;
            }
        }
        case actl_data: {
            analyzer_mst.valid <= 1;
            analyzer_mst.data <= apb_state.control.data[4;0];
            apb_state.control.data <= apb_state.control.data>>4;
            apb_state.control.nybbles <= apb_state.control.nybbles-1;
            if (apb_state.control.nybbles==0) {
                analyzer_mst.valid <= 0;
                analyzer_mst.data <= 0;
                apb_state.control.state <= actl_idle;
                apb_state.control.write_data <= 0;
            }
        }            
        }
        if (apb_state.access==access_write_mux_control) {
            apb_state.control.enable        <= apb_request.pwdata[0];
            apb_state.control.write_data    <= apb_request.pwdata[1];
            apb_state.control.nybbles       <= apb_request.pwdata[3;4];
            apb_state.control.data          <= apb_request.pwdata[24;8];
        }            
    }

    /*b APB interface
     */
    apb_interface "APB interface": {
        /*b Handle APB read data - may affect pready */
        apb_read_trace      = 0;
        apb_response = {*=0, pready=1};
        part_switch (apb_state.access) {
        case access_read_status: {
            apb_response.prdata[0] = apb_trigger_reset;
            apb_response.prdata[1] = apb_trigger_enable;
            apb_response.prdata[2] = apb_trace_readback;
            apb_response.prdata[3] = apb_trace_valid; // note not stable - need to fix
            apb_response.prdata[4] = trigger_reset;   // note not stable - need to fix
            apb_response.prdata[5] = trigger_enable;  // note not stable - need to fix
            apb_response.prdata[6] = trigger_done;    // note not stable - need to fix
            apb_response.prdata[7] = trigger_circular;
            apb_response.prdata[8] = analyzer_tgt_r.enable_return;
            apb_response.prdata[9] = analyzer_tgt_r.selected;
            apb_response.prdata[2;10] = trigger_stage;  // note not stable - need to fix
            apb_response.prdata[analyzer_trigger_counter_width;16] = trigger_residence;  // note not stable - need to fix
        }
        case access_read_trace_data: {
            apb_response.prdata = apb_trace_data;
            apb_read_trace      = 1;
        }
        }

        /*b Handle APB writes - may affect pready */
        part_switch (apb_state.access) {
        case access_write_config: {
            apb_trigger_reset  <= apb_request.pwdata[0];
            apb_trigger_enable <= apb_request.pwdata[1];
            apb_trace_readback <= apb_request.pwdata[2];
            trigger_circular   <= apb_request.pwdata[7];
            apb_trigger_stage  <= apb_request.pwdata[analyzer_trigger_depth_log;8];
        }
        case access_write_trigger: {
            trigger[ apb_trigger_stage ] <= { counter=apb_request.pwdata[analyzer_trigger_counter_width;0],
                    if_true=apb_request.pwdata[analyzer_trigger_depth_log;16],
                    action_if_true=apb_request.pwdata[3;20],
                    if_false=apb_request.pwdata[analyzer_trigger_depth_log;24],
                    action_if_false=apb_request.pwdata[3;28] };
        }
        case access_write_mask: {
            trigger[ apb_trigger_stage ].mask <= apb_request.pwdata[ analyzer_trigger_signal_width; 0];
        }
        case access_write_compare: {
            trigger[ apb_trigger_stage ].compare <= apb_request.pwdata[ analyzer_trigger_signal_width; 0];
        }
        }

        /*b Decode access */
        apb_state.access <= access_none;
        part_switch (apb_request.paddr[4;0]) {
        case apb_address_config_byte_0: {
            apb_state.access <= apb_request.pwrite ? access_write_config_byte_0 : access_none;
        }
        case apb_address_config_byte_1: {
            apb_state.access <= apb_request.pwrite ? access_write_config_byte_1 : access_none;
        }
        case apb_address_config_byte_2: {
            apb_state.access <= apb_request.pwrite ? access_write_config_byte_2 : access_none;
        }
        case apb_address_config_byte_3: {
            apb_state.access <= apb_request.pwrite ? access_write_config_byte_3 : access_none;
        }
        case apb_address_action_source_0: {
            apb_state.access <= apb_request.pwrite ? access_write_action_source_0 : access_none;
        }
        case apb_address_action_source_1: {
            apb_state.access <= apb_request.pwrite ? access_write_action_source_1 : access_none;
        }
        case apb_address_cfg: {
            apb_state.access <= apb_request.pwrite ? access_write_config : access_none;
        }
        case apb_address_trace_data: {
            apb_state.access <= apb_request.pwrite ? access_none : access_read_trace_data;
        }
        }
        if (!apb_request.psel || (apb_request.penable && apb_response.pready)) {
            apb_state.access <= access_none;
        }

    }

    /*b Done
     */
}
