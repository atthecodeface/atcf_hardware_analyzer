/*a Includes
 */
include "analyzer.h"
include "analyzer_trigger.h"
include "clocking::clock_timer.h"
include "std::valid_data.h"

/*a Types
 */
/*t t_timer_combs
 */
typedef struct
{
    bit[32] value;
    bit[32] timer_delta;
} t_timer_combs;

/*t t_timer_state
 */
typedef struct
{
    bit[32] value;
    t_vdata_32 recorded_value;
    bit[32] timer_delta "Valid if recorded_value is valid";
} t_timer_state;

/*a Module
 */
module analyzer_trigger_timer( clock clk,
                               input bit reset_n,

                               input  t_analyzer_trigger_cfg trigger_cfg,
                               input  t_analyzer_trigger_ctl trigger_ctl,
                               input t_timer_value timer_value,
                               input bit record_time,
                               output t_analyzer_trigger_timer trigger_timer
    )
"""
This module is designed to trigger on an 8-bit mask/match of one byte of the input data

The output data can be data in or the timer value
"""

{
    /*b Default clock and reset
     */
    default clock clk;
    default reset active_low reset_n;

    /*b State and combs */
    clocked t_timer_state timer_state = {*=0};
    comb t_timer_combs timer_combs;

    /*b Timer value outputs
     */
    timer_value_outputs "Timer value outputs logic": {
        trigger_timer.value = timer_state.value;
        trigger_timer.timer_delta = timer_combs.timer_delta;
        trigger_timer.recorded_value = timer_state.recorded_value;
        trigger_timer.recorded_delta.valid = timer_state.recorded_value.valid;
        trigger_timer.recorded_delta.data = timer_state.timer_delta;
    }

    /*b Timer value state
     */
    timer_value_logic "Timer value logic": {
        timer_combs.value = timer_value.value[32;0];
        full_switch (trigger_cfg.timer_div) {
        case 2b00: {
            timer_combs.value = timer_value.value[32;0];
        }
        case 2b01: {
            timer_combs.value = timer_value.value[32;8];
        }
        case 2b10: {
            timer_combs.value = timer_value.value[32;16];
        }
        case 2b11: {
            timer_combs.value = timer_state.value+1;
        }
        }

        timer_state.value <= timer_combs.value;
        timer_combs.timer_delta = timer_state.value - timer_state.recorded_value.data;
        if (timer_state.recorded_value.valid) {
            timer_state.timer_delta <= timer_combs.timer_delta;
        }

        if (record_time) {
            timer_state.recorded_value.valid <= 1;
            timer_state.recorded_value.data <= timer_state.value;
            timer_state.timer_delta <= 0;
        }

        if (trigger_ctl.clear) {
            timer_state <= {*=0};
        }

        if (!trigger_ctl.enable) {
            timer_state <= timer_state;
        }

    }
}
