/*a Includes
 */
include "analyzer.h"

/*a Types */
/*t t_actl_fsm_state
 */
typedef fsm {
    actl_fsm_idle;
    actl_fsm_select_at;
    actl_fsm_select_run_all;
    actl_fsm_select_run_clear_enable;
    actl_fsm_write_data;
    actl_fsm_completed;
} t_actl_fsm_state;

/*t t_actl_state */
typedef struct {
    t_actl_fsm_state fsm_state;
    t_analyzer_mst mst;
    t_analyzer_tgt tgt;
    bit[60] data;
    bit[4] count;
    bit completed;
} t_actl_state;

/*a Module
 */
module analyzer_control_master( clock clk,
                                input bit reset_n,

                                input t_analyzer_mst_ctl mst_ctl,
                                output t_analyzer_mst_ctl_resp mst_ctl_resp,

                                output  t_analyzer_mst  analyzer_mst,
                                input t_analyzer_tgt  analyzer_tgt "Data not used"

    )
"""
This module drives the analyzer_mst bus as the root of the control bus.

A select transaction with data of 'count' drives enable down the
analyzer control chain and waits for it to return high; it sets
'select' high (and keeps it there) after 'count' cycles; this is used
to select a particular target on the chain.

A select write with data 0 selects *no* targets; it clears select and
then drives enable high, and waits (counting) until enable_return is
high. The count, at this point, indicates the length of the chain. A
select write with data 1 does the same by keeping the select signal
high for this duration.

[ Why would one do a select with data of 1? ]

A select write with top data bit set forces enable to be clear, and it
waits until enable_return is clear, counting.

Once a select has completed, data can be written to the selected
target by a 'write data' command; this shifts data in from the bottom,
reversing the nybbles; nybbles are shifted out as they are written,
and data stops being written when it is zero - so the last nybble that
is to be written (the bottom nybble of data at the target) must be
non-zero. Note that if a target is configured with a trace width of
less than four 32-bit values then it will include a multiplexer
selected by the last nybble written.

Usage

Perform a select write with data 0, to count the length of the
analyzer control chain; when the status read has top bit set the count
will be correct. This clears the drivers as well as counting.

Clear the enable with a select write with data with the top bit set;
wait for that to complete.

Select a specific target by first clearing the enable, then performing
a 'select_at'.

"""

{
    /*b Default clock and reset
     */
    default clock clk;
    default reset active_low reset_n;

    /*b Internal state
     */
    clocked t_actl_state actl_state = {*=0};

    /*b Capture analyzer_tgt bus
     */
    analyzer_tgt_capture "Record analyzer_tgt": {
        mst_ctl_resp = {
            completed = actl_state.completed,
            selected = actl_state.tgt.selected,
            count = actl_state.data[16;0]
        };
        if (actl_state.mst.enable ||
            actl_state.mst.select ||
            actl_state.tgt.enable_return ||
            analyzer_tgt.enable_return) {
            actl_state.tgt <= analyzer_tgt;
        }
    }
        
    /*b Analyzer control FSM
     */
    analyzer_control_fsm "Analyzer control FSM logic": {
        full_switch (actl_state.fsm_state) {
        case actl_fsm_idle: {
            if (mst_ctl.actl_op != actl_op_none) {
                actl_state.completed <= 0;
                actl_state.mst <= {*=0};
                actl_state.data <= 0;
            }
            full_switch (mst_ctl.actl_op) {
            case actl_op_select: {
                actl_state.fsm_state <= actl_fsm_select_at;
                actl_state.data[32;0] <= mst_ctl.data[32;0];
            }
            case actl_op_clear_enable: {
                actl_state.fsm_state <= actl_fsm_select_run_clear_enable;
            }
            case actl_op_select_all: {
                actl_state.fsm_state <= actl_fsm_select_run_all;
                actl_state.mst.select <= 1;
            }
            case actl_op_select_none: {
                actl_state.fsm_state <= actl_fsm_select_run_all;
            }
            case actl_op_write_data: {
                actl_state.fsm_state <= actl_fsm_write_data;
                actl_state.mst <= actl_state.mst;
                actl_state.mst.valid <= 1;
                actl_state.mst.data <= mst_ctl.data[4;60];
                actl_state.data <= mst_ctl.data[60; 0];
                actl_state.count <= 15;
            }
        }
        }
        case actl_fsm_select_run_all: {
            actl_state.mst.enable <= 1;
            if (actl_state.tgt.enable_return) {
                actl_state.fsm_state <= actl_fsm_completed;
            }
            actl_state.data[32;0] <= actl_state.data[32;0] + 1;
        }
        case actl_fsm_select_run_clear_enable: {
            if (!actl_state.tgt.enable_return) {
                actl_state.fsm_state <= actl_fsm_completed;
            }
            actl_state.data[32;0] <= actl_state.data[32;0] + 1;
        }
        case actl_fsm_select_at: {
            actl_state.mst.enable <= 1;
            actl_state.mst.select <= 0;
            if (actl_state.data[32;0] == 0) {
                actl_state.mst.select <= 1;
            }
            if (actl_state.tgt.enable_return) {
                actl_state.fsm_state <= actl_fsm_completed;
            }
            actl_state.data[32;0] <= actl_state.data[32;0] - 1;
        }
        case actl_fsm_write_data: {
            actl_state.mst.valid <= 1;
            actl_state.mst.data <= actl_state.data[4;56];
            actl_state.data <= actl_state.data << 4;
            if (actl_state.count == 0) {
                actl_state.fsm_state <= actl_fsm_completed;
                actl_state.mst.valid <= 0;
            }
            actl_state.count <= actl_state.count-1;
        }
        case actl_fsm_completed: {
            actl_state.fsm_state <= actl_fsm_idle;
            actl_state.completed <= 1;
        }
        }            

        analyzer_mst = actl_state.mst;
    }

    /*b Done
     */
}
