/*a Includes
 */
include "apb::apb.h"
include "analyzer.h"
include "analyzer_modules.h"
include "std::srams.h"

/*a Constants */
constant integer apb_reads = 0;

/*a Types */
/*t t_apb_address
 * APB address map, used to decode paddr
 *
 * The APB decodes to trace/trigger/filter, then which of those, and then which fields
 *
 * Could add timer as an optional 4th
 */
typedef enum [4] {
    apb_address_filter  = 0,
    apb_address_trigger = 1,
    apb_address_trace   = 2,
} t_apb_address_kind;

/*t t_apb_address_trace
 * APB address map for trace
 *
 *
 */
typedef enum [4] {
    apb_trace_base               = 0,
    apb_trace_fifos              = 1,
    apb_trace_offset_base        = 2,
    apb_trace_offset_shift_size  = 3,
    apb_trace_value_0_base       = 4,
    apb_trace_value_0_shift_size = 5,
    apb_trace_value_1_base       = 6,
    apb_trace_value_1_shift_size = 7,
} t_apb_trace_ofs;

/*t t_apb_address_trigger
 * APB address map for trigger
 *
 *
 */
typedef enum [4] {
    apb_trigger_base               = 0,
    apb_trigger_match_data_src     = 1, // 12
    apb_trigger_match_byte_0          = 4, // 22
    apb_trigger_match_byte_1          = 5, // 22
    apb_trigger_match_byte_2          = 6, // 22
    apb_trigger_match_byte_3          = 7, // 22
    apb_trigger_set_0    = 8, // 24 - map 4-bit bundle of matches to one of 8 sets-of-actions
    apb_trigger_set_1    = 9, // 24 - map 4-bit bundle of matches to one of 8 sets-of-actions
    apb_trigger_actions_0       = 10, // 4 * 6 - four sets-of-actions
    apb_trigger_actions_1       = 11, // 4 * 6 - four sets-of-actions
} t_apb_trigger_ofs;

/*t t_apb_address_filter
 * APB address map for filter
 *
 *
 */
typedef enum [4] {
    apb_filter_base       = 0,
    apb_filter_mask_0     = 8,
    apb_filter_mask_1     = 9,
    apb_filter_mask_2     = 10,
    apb_filter_mask_3     = 11,
    apb_filter_value_0    = 12,
    apb_filter_value_1    = 13,
    apb_filter_value_2    = 14,
    apb_filter_value_3    = 15,
} t_apb_filter_ofs;

/*t t_access
 * APB access that is in progress; a decode of psel and paddr
 */
typedef enum [3] {
    access_none        "No access being performed",
    access_write_trigger  "Write data to trigger cfg",
    access_write_trace    "Write data to trace cfg",
    access_write_filter   "Write data to filter cfg",
    access_read_trigger  "Read data from trigger cfg",
    access_read_trace    "Read data from trace cfg",
    access_read_filter   "Read data from filter cfg",
} t_access;

/*t t_apb_combs */
typedef struct {
    bit[32] trigger_read_data;
    bit[32] trace_read_data;
    bit[32] filter_read_data;
} t_apb_combs;

/*t t_apb_state */
typedef struct {
    t_access access;
    bit[32] write_data;
    bit[4] ofs;
    t_analyzer_filter_cfg filter_cfg;
    t_analyzer_trigger_cfg trigger_cfg;
    t_analyzer_trace_cfg trace_cfg;
} t_apb_state;

/*a Module
 */
module apb_target_analyzer_cfg( clock clk,
                                input bit reset_n,

                                input  t_apb_request  apb_request  "APB request",
                                output t_apb_response apb_response "APB response",

                                output  t_analyzer_filter_cfg filter_cfg,
                                output  t_analyzer_trigger_cfg trigger_cfg,
                                output  t_analyzer_trace_cfg trace_cfg
    )
"""
This module provides configuration for logic analyzers from APB.

Most of the configuration can be configured to be write-only; this is
because the analyzer is designed to be purely used for silicon debug,
and is not really expected to be exposed to most software, let alone
'consumers'.

This also enables designs that do not use some of the configuration to
synthesize out the unused configuration flops.
                                                                  
"""

{
    /*b Default clock and reset
     */
    default clock clk;
    default reset active_low reset_n;

    /*b APB state and combs
     */
    clocked t_apb_state apb_state = {*=0};
    comb t_apb_combs apb_combs;

    /*b Drive the output configuration
     */
    drive_outputs "Drive the ouputs": {
        filter_cfg = apb_state.filter_cfg;
        trigger_cfg = apb_state.trigger_cfg;
        trace_cfg = apb_state.trace_cfg;
    }

    /*b APB read
     */
    apb_reads "APB reads": {

        /*b Handle APB read data - may affect pready */
        apb_response = {*=0, pready=1};
        part_switch (apb_state.access) {
        case access_read_trigger: {
            apb_response.prdata |= apb_combs.trigger_read_data;
        }
        case access_read_filter: {
            apb_response.prdata |= apb_combs.filter_read_data;
        }
        case access_read_trace: {
            apb_response.prdata |= apb_combs.trace_read_data;
        }
        }
    }
    
    /*b APB interface state
     */
    apb_interface "APB interface": {

        /*b Decode access */
        apb_state.access <= access_none;
        apb_state.ofs <= apb_request.paddr[4;0];
        apb_state.write_data <= apb_request.pwdata;
        part_switch (apb_request.paddr[4;4]) {
        case apb_address_trigger: {
            apb_state.access <= apb_request.pwrite ? access_write_trigger: access_read_trigger;
        }
        case apb_address_trace: {
            apb_state.access <= apb_request.pwrite ? access_write_trace: access_read_trace;
        }
        case apb_address_filter: {
            apb_state.access <= apb_request.pwrite ? access_write_filter: access_read_filter;
        }
        }
        if (!apb_request.psel || (apb_request.penable && apb_response.pready)) {
            apb_state.access <= access_none;
            apb_state.ofs <= apb_state.ofs;
            apb_state.write_data <= apb_state.write_data;
        }
    }

    /*b Filter config
     */
    filter_config_logic "Filter configuration logic": {
        apb_state.trace_cfg <= apb_state.trace_cfg;

        /*b Keep state */
        full_switch (apb_state.ofs) {
        case apb_filter_base: {
            apb_state.filter_cfg.enable <= apb_state.write_data[0];
            apb_state.filter_cfg.accept_unchanging <= apb_state.write_data[1];
        }
        case apb_filter_mask_0: {
            apb_state.filter_cfg.mask.data_0 <= apb_state.write_data;
        }
        case apb_filter_mask_1: {
            apb_state.filter_cfg.mask.data_1 <= apb_state.write_data;
        }
        case apb_filter_mask_2: {
            apb_state.filter_cfg.mask.data_2 <= apb_state.write_data;
        }
        case apb_filter_mask_3: {
            apb_state.filter_cfg.mask.data_3 <= apb_state.write_data;
        }
        case apb_filter_value_0: {
            apb_state.filter_cfg.value.data_0 <= apb_state.write_data;
        }
        case apb_filter_value_1: {
            apb_state.filter_cfg.value.data_1 <= apb_state.write_data;
        }
        case apb_filter_value_2: {
            apb_state.filter_cfg.value.data_2 <= apb_state.write_data;
        }
        case apb_filter_value_3: {
            apb_state.filter_cfg.value.data_3 <= apb_state.write_data;
        }
        }

        full_switch (apb_state.ofs) {
        case apb_trigger_base: {
            apb_state.trigger_cfg.enable <= apb_state.write_data[0];
            apb_state.trigger_cfg.clear <= apb_state.write_data[1];
            apb_state.trigger_cfg.start <= apb_state.write_data[2];
            apb_state.trigger_cfg.stop <= apb_state.write_data[3];
            apb_state.trigger_cfg.timer_div <= apb_state.write_data[2; 8];
        }
        case apb_trigger_match_data_src: {
            apb_state.trigger_cfg.data_src_0 <= apb_state.write_data[2; 0];
            apb_state.trigger_cfg.data_src_1 <= apb_state.write_data[2; 8];
            apb_state.trigger_cfg.match_data_src_0 <= apb_state.write_data[3; 16];
            apb_state.trigger_cfg.match_data_src_1 <= apb_state.write_data[3; 24];
        }
        case apb_trigger_match_byte_0: {
            apb_state.trigger_cfg.tb_0.ignore_valid <= apb_state.write_data[0];
            apb_state.trigger_cfg.tb_0.byte_sel <= apb_state.write_data[3; 8];
            apb_state.trigger_cfg.tb_0.cond_sel <= apb_state.write_data[2; 12];
            apb_state.trigger_cfg.tb_0.mask <= apb_state.write_data[8; 16];
            apb_state.trigger_cfg.tb_0.match <= apb_state.write_data[8; 24];
        }
        case apb_trigger_match_byte_1: {
            apb_state.trigger_cfg.tb_1.ignore_valid <= apb_state.write_data[0];
            apb_state.trigger_cfg.tb_1.byte_sel <= apb_state.write_data[3; 8];
            apb_state.trigger_cfg.tb_1.cond_sel <= apb_state.write_data[2; 12];
            apb_state.trigger_cfg.tb_1.mask <= apb_state.write_data[8; 16];
            apb_state.trigger_cfg.tb_1.match <= apb_state.write_data[8; 24];
        }
        case apb_trigger_match_byte_2: {
            apb_state.trigger_cfg.tb_2.ignore_valid <= apb_state.write_data[0];
            apb_state.trigger_cfg.tb_2.byte_sel <= apb_state.write_data[3; 8];
            apb_state.trigger_cfg.tb_2.cond_sel <= apb_state.write_data[2; 12];
            apb_state.trigger_cfg.tb_2.mask <= apb_state.write_data[8; 16];
            apb_state.trigger_cfg.tb_2.match <= apb_state.write_data[8; 24];
        }
        case apb_trigger_match_byte_3: {
            apb_state.trigger_cfg.tb_3.ignore_valid <= apb_state.write_data[0];
            apb_state.trigger_cfg.tb_3.byte_sel <= apb_state.write_data[3; 8];
            apb_state.trigger_cfg.tb_3.cond_sel <= apb_state.write_data[2; 12];
            apb_state.trigger_cfg.tb_3.mask <= apb_state.write_data[8; 16];
            apb_state.trigger_cfg.tb_3.match <= apb_state.write_data[8; 24];
        }
        case apb_trigger_set_0: {
            apb_state.trigger_cfg.action_set[24; 0] <= apb_state.write_data[24; 0];
        }
        case apb_trigger_set_1: {
            apb_state.trigger_cfg.action_set[24; 24] <= apb_state.write_data[24; 0];
        }
        case apb_trigger_actions_0: {
            apb_state.trigger_cfg.actions_0.halt_capture       <= apb_state.write_data[0];
            apb_state.trigger_cfg.actions_0.record_data        <= apb_state.write_data[1];
            apb_state.trigger_cfg.actions_0.record_time        <= apb_state.write_data[2];
            apb_state.trigger_cfg.actions_0.record_invalidate  <= apb_state.write_data[3];
            apb_state.trigger_cfg.actions_0.capture_data       <= apb_state.write_data[2; 4];

            apb_state.trigger_cfg.actions_1.halt_capture       <= apb_state.write_data[8];
            apb_state.trigger_cfg.actions_1.record_data        <= apb_state.write_data[9];
            apb_state.trigger_cfg.actions_1.record_time        <= apb_state.write_data[10];
            apb_state.trigger_cfg.actions_1.record_invalidate  <= apb_state.write_data[11];
            apb_state.trigger_cfg.actions_1.capture_data       <= apb_state.write_data[2; 12];

            apb_state.trigger_cfg.actions_2.halt_capture       <= apb_state.write_data[16];
            apb_state.trigger_cfg.actions_2.record_data        <= apb_state.write_data[17];
            apb_state.trigger_cfg.actions_2.record_time        <= apb_state.write_data[18];
            apb_state.trigger_cfg.actions_2.record_invalidate  <= apb_state.write_data[19];
            apb_state.trigger_cfg.actions_2.capture_data       <= apb_state.write_data[2; 20];

            apb_state.trigger_cfg.actions_3.halt_capture       <= apb_state.write_data[24];
            apb_state.trigger_cfg.actions_3.record_data        <= apb_state.write_data[25];
            apb_state.trigger_cfg.actions_3.record_time        <= apb_state.write_data[26];
            apb_state.trigger_cfg.actions_3.record_invalidate  <= apb_state.write_data[27];
            apb_state.trigger_cfg.actions_3.capture_data       <= apb_state.write_data[2; 28];
        }
        case apb_trigger_actions_1: {
            apb_state.trigger_cfg.actions_4.halt_capture       <= apb_state.write_data[0];
            apb_state.trigger_cfg.actions_4.record_data        <= apb_state.write_data[1];
            apb_state.trigger_cfg.actions_4.record_time        <= apb_state.write_data[2];
            apb_state.trigger_cfg.actions_4.record_invalidate  <= apb_state.write_data[3];
            apb_state.trigger_cfg.actions_4.capture_data       <= apb_state.write_data[2; 4];

            apb_state.trigger_cfg.actions_5.halt_capture       <= apb_state.write_data[8];
            apb_state.trigger_cfg.actions_5.record_data        <= apb_state.write_data[9];
            apb_state.trigger_cfg.actions_5.record_time        <= apb_state.write_data[10];
            apb_state.trigger_cfg.actions_5.record_invalidate  <= apb_state.write_data[11];
            apb_state.trigger_cfg.actions_5.capture_data       <= apb_state.write_data[2; 12];

            apb_state.trigger_cfg.actions_6.halt_capture       <= apb_state.write_data[16];
            apb_state.trigger_cfg.actions_6.record_data        <= apb_state.write_data[17];
            apb_state.trigger_cfg.actions_6.record_time        <= apb_state.write_data[18];
            apb_state.trigger_cfg.actions_6.record_invalidate  <= apb_state.write_data[19];
            apb_state.trigger_cfg.actions_6.capture_data       <= apb_state.write_data[2; 20];

            apb_state.trigger_cfg.actions_7.halt_capture       <= apb_state.write_data[24];
            apb_state.trigger_cfg.actions_7.record_data        <= apb_state.write_data[25];
            apb_state.trigger_cfg.actions_7.record_time        <= apb_state.write_data[26];
            apb_state.trigger_cfg.actions_7.record_invalidate  <= apb_state.write_data[27];
            apb_state.trigger_cfg.actions_7.capture_data       <= apb_state.write_data[2; 28];
        }
        default: {
            apb_state.trigger_cfg <= apb_state.trigger_cfg;
        }
        }
        if (apb_state.access != access_write_filter) {
            apb_state.filter_cfg <= apb_state.filter_cfg;
        }
        if (apb_state.access != access_write_trigger) {
            apb_state.trigger_cfg <= apb_state.trigger_cfg;
        }

        apb_combs.trigger_read_data = 0;
        apb_combs.trace_read_data = 0;
        apb_combs.filter_read_data = 0;
        if (!(apb_reads&1)) {
            apb_combs.filter_read_data = 0;
        }
        if (!(apb_reads&2)) {
            apb_combs.trigger_read_data = 0;
        }
        if (!(apb_reads&4)) {
            apb_combs.trace_read_data = 0;
        }

    }

    /*b Done
     */
}
