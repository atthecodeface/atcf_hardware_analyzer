/** @copyright (C) 2020,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   analyzer_target.cdl
 * @brief  Standard target for the analyzer bus
 *

 */

/*a Includes
 */
include "analyzer.h"
include "std::tech_sync.h"

/*a Types
*/
/*t t_out_combs */
typedef struct {
    bit[4] toggle_difference;
} t_out_combs;

/*t t_out_state */
typedef struct {
    bit[2] next_data_out;
    bit[4] toggle;
    t_analyzer_data data_out;
} t_out_state;

/*t t_in_state */
typedef struct {
    bit[2] next_data_in;
    bit[4] valid_toggle;
} t_in_state;

/*a Module
 */
/*m analyzer_async_data_slow_to_fast
 *
 * Analyzer data clock domain crossing
 *
 */
module analyzer_async_data_slow_to_fast( clock clk_in,
                                         clock clk_out,
                                         input bit reset_n,

                                         input t_analyzer_data analyzer_data_in,
                                         output t_analyzer_data analyzer_data_out
    )
{
    /*b Clock in state */
    default clock clk_in;
    default reset active_low reset_n;
    clocked t_in_state         in_state = {*=0};
    clocked t_analyzer_data[4] data_buffer  = {*=0};

    /*b Clock out state */
    default clock clk_out;
    default reset active_low reset_n;
    comb    t_out_combs        out_combs;
    clocked t_out_state        out_state = {*=0};
    net bit[4] out_valid_toggle;

    /*b Clock in logic */
    clock_in_logic : {
        if (analyzer_data_in.valid) {
            in_state.valid_toggle[in_state.next_data_in] <= !in_state.valid_toggle[in_state.next_data_in];
            data_buffer[in_state.next_data_in].valid <= 0;
            data_buffer[in_state.next_data_in].data  <= analyzer_data_in.data;
            in_state.next_data_in <= in_state.next_data_in + 1;
        }
    }        
        
    /*b Clock out logic */
    clock_out_logic : {
        
        for (i; 4) {
            tech_sync_bit toggle_sync_flops[i](clk <- clk_out, reset_n <= reset_n,
                                               d <= in_state.valid_toggle[i],
                                               q => out_valid_toggle[i] );
        }
        out_combs.toggle_difference = out_valid_toggle ^ out_state.toggle;

        out_state.data_out.valid <= 0;
        if (out_combs.toggle_difference[out_state.next_data_out]) {
            out_state.data_out.valid                  <= 1;
            out_state.data_out.data                   <= data_buffer[out_state.next_data_out].data;
            out_state.toggle[out_state.next_data_out] <= !out_state.toggle[out_state.next_data_out];
            out_state.next_data_out <= out_state.next_data_out + 1;
        }
        analyzer_data_out = out_state.data_out;
        /*b All done */
    }

    /*b All done */
}
