/*a Includes */
include "apb::apb.h"
include "apb::apb_masters.h"
include "std::srams.h"
include "utils::fifo_status.h"
include "utils::debug.h"
include "utils::debug_modules.h"
include "clocking::clock_timer.h"
include "clocking::clock_timer_modules.h"

include "analyzer.h"
include "analyzer_modules.h"
include "tb_analyzer_modules.h"

/*a Module */
module tb_analyzer_dbg( clock clk,
                        input bit reset_n,

                        input t_dbg_master_request dbg_master_req,
                        output t_dbg_master_response dbg_master_resp
)
{

    /*b Nets */
    default clock clk;
    default reset active_low reset_n;
    net t_dbg_master_response dbg_master_resp;

    net t_dbg_master_request  dbg_master_req_fifo;
    net t_dbg_master_request  dbg_master_req_apb;
    net t_dbg_master_response dbg_master_resp_fifo;
    net t_dbg_master_response dbg_master_resp_apb;

    net t_analyzer_mst analyzer_mst;
    net t_analyzer_tgt analyzer_tgt;
    net t_analyzer_trace_op4 analyzer_trace_op;

    default clock clk;
    default reset active_low reset_n;

    net  t_analyzer_data4 analyzer_data_filtered;
    net  t_analyzer_data4 analyzer_data_triggered;

    net  t_analyzer_filter_cfg filter_cfg;
    net  t_analyzer_trigger_cfg trigger_cfg;
    net  t_analyzer_trace_cfg trace_cfg;
    comb  t_timer_control_full timer_ctl;
    net t_timer_value  timer_value;
    
    net t_fifo_status[2] trace_fifo_status;

    comb t_analyzer_trace_access_req trace_access_req;
    comb bit[4] trace_access_valid;
    net t_analyzer_trace_access_resp trace_access_resp;
    net bit trace_access_rdy;

    net t_apb_request             apb_request;
    comb t_apb_response            apb_response;

    comb  t_apb_request  apb_request_ctl  "APB request to target ctl";
    comb  t_apb_request  apb_request_cfg  "APB request to target cfg";
    comb  t_apb_request  apb_request_src  "APB request to target src";
    net t_apb_response apb_response_ctl "APB response from target ctl";
    net t_apb_response apb_response_cfg "APB response from target cfg";
    net t_apb_response apb_response_src "APB response from target src";

    comb t_dbg_master_response resp_none;
    net bit dbg_pop_fifo;

    /*b Instantiations */
    instantiations: {
        apb_response = {*=0};
        apb_response |= apb_response_cfg;
        apb_response |= apb_response_ctl;
        apb_response |= apb_response_src;

        apb_response.pready = (apb_response_cfg.pready &
                               apb_response_ctl.pready &
                               apb_response_src.pready);

        apb_request_cfg = apb_request;
        apb_request_ctl = apb_request;
        apb_request_src = apb_request;
        apb_request_cfg.psel = apb_request.psel && (apb_request.paddr[2;10] == 2b00);
        apb_request_ctl.psel = apb_request.psel && (apb_request.paddr[2;10] == 2b01);
        apb_request_src.psel = apb_request.psel && (apb_request.paddr[2;10] == 2b11);

        timer_ctl = {*=0};

        trace_access_req = {*=0};
        trace_access_req.read_enable = 1;
        trace_access_req.id = 2b11;
        trace_access_req.address_op = atr_address_op_pop;

        trace_access_valid = 0;
        trace_access_valid[0] = dbg_pop_fifo;

        resp_none = {*=0};
        
        dbg_master_mux mux( clk <- clk,
                                 reset_n <= reset_n,
                                 dbg_master_req <= dbg_master_req,
                                 dbg_master_resp => dbg_master_resp,
                                 req1 => dbg_master_req_fifo,
                                 req2 => dbg_master_req_apb,
                                 resp0 <= resp_none,
                                 resp1 <= dbg_master_resp_fifo,
                                 resp2 <= dbg_master_resp_apb,
                                 resp3 <= resp_none
            );

        dbg_master_fifo_sink dut( clk <- clk,
                                 reset_n <= reset_n,
                                  dbg_master_req <= dbg_master_req_fifo,
                                  dbg_master_resp => dbg_master_resp_fifo,
                                  fifo_status <= trace_fifo_status[0],
                                  data0 <= bundle(32b0, trace_access_resp.data),
                                  data1 <= 0,
                                  data2 <= 0,
                                  data3 <= 0,
                                  pop_rdy <= trace_access_rdy,
                                  data_valid <= trace_access_resp.valid && (trace_access_resp.id==2b11),
                                  pop_fifo => dbg_pop_fifo
            );

        apb_script_master apb( clk <- clk,
                       reset_n <= reset_n,

                       dbg_master_req <= dbg_master_req_apb,
                       dbg_master_resp => dbg_master_resp_apb,
                       apb_request => apb_request,
                       apb_response  <= apb_response );


        apb_target_analyzer_ctl ctl( clk <- clk,
                                     reset_n <= reset_n,
                                     apb_request <= apb_request_ctl,
                                     apb_response => apb_response_ctl,
                                     analyzer_mst => analyzer_mst,
                                     analyzer_tgt <= analyzer_tgt
            );

        apb_target_analyzer_cfg cfg( clk <- clk,
                                     reset_n <= reset_n,
                                     apb_request <= apb_request_cfg,
                                     apb_response => apb_response_cfg,
                                     filter_cfg => filter_cfg,
                                     trigger_cfg => trigger_cfg,
                                     trace_cfg => trace_cfg );

        clock_timer clk_timer( clk<-clk, reset_n<=reset_n,
                               timer_control <= timer_ctl,
                               timer_value => timer_value);

        tb_apb_target_analyzer_src src( clk <- clk, reset_n <= reset_n,
                                     apb_request <= apb_request_src,
                                     apb_response => apb_response_src,
                             analyzer_mst <= analyzer_mst,
                             analyzer_tgt => analyzer_tgt
            );

        analyzer_trace_filter filter( clk <- clk, reset_n <= reset_n,
                                      din <= analyzer_tgt.data,
                                      dout => analyzer_data_filtered,
                                      filter_cfg <= filter_cfg );

        analyzer_trigger_simple trigger(  clk <- clk, reset_n <= reset_n,
                                          din <= analyzer_data_filtered,
                                          dout => analyzer_data_triggered,
                                          trace_op => analyzer_trace_op,
                                          timer_value <= timer_value,
                                          trigger_cfg_in <= trigger_cfg );

        analyzer_trace_ram trace(  clk <- clk, reset_n <= reset_n,
                                   trace_op <= analyzer_trace_op,
                                   din <= analyzer_data_triggered,
                                   fifo_status_l => trace_fifo_status[0],
                                   fifo_status_h => trace_fifo_status[1],

                                   trace_access_req <= trace_access_req,
                                   trace_access_rdy => trace_access_rdy,
                                   trace_access_valid <= trace_access_valid[2;0],
                                   trace_access_resp => trace_access_resp,

                                   trace_cfg <= trace_cfg );

    }
}
