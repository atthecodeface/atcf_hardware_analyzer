/*a Includes
 */
include "analyzer.h"
include "analyzer_modules.h"
include "analyzer_trace_ram.h"
include "utils::fifo_status.h"
include "clocking::clock_timer.h"
include "std::srams.h"

/*a Types */
/*t t_timer_state
 */
typedef struct
{
    bit[32] value;
} t_timer_state;

/*t t_recorded_state
 */
typedef struct
{
    bit[32] timer;
    bit[32][2] data;
} t_recorded_state;

/*t t_match_combs
 */
typedef struct
{
    t_analyzer_data4 data;
    bit data_changing;
    bit[2] matched;
    bit record_data;
    bit record_time;
    bit[2] capture_data;
} t_match_combs;

/*a Module
 */
module analyzer_trigger_simple( clock clk,
                           input bit reset_n,

                           input  t_analyzer_data4  din,
                           output  t_analyzer_data4 dout,

                           output  t_analyzer_trace_op4 trace_op,
                           input t_timer_value timer_value,

                           input  t_analyzer_trigger_cfg trigger_cfg
 )
"""

For each byte mask match of N:

* Select which din

* Select byte of data

* One mask/match per selected byte yields 'match' and 'match changed' (6 conditions in fact)

Yields 6*N bits

Combining 6*N bits:

* Two cfgs of select-bit-of-6 for each N byte mask match, plus 'only if any data changing'

* cfg has independent action options of record time; record data; capture data out 0; capture data out 1

* output can be configured to be time, time delta, data, data delta.


So some configurations:


* Record time that state machine is not idle; captures time leaves idle, time enters idle, and deltas

* byte mask/match 0 on din.data0[8;0] == 8b_xxx000xx (idle state of fsm)

* If BMM 0 set: record time

* If BMM 0 set and changed: capture dout_0 = time delta, capture dout_1 = time value


* Record FSM state and time since last idle.

* byte mask/match 0 on din.data0[8;0] == 8b_xxx000xx (idle state of fsm)

* byte mask/match 1 on din.data0[8;0] == 8b_xxxSSSxx (other state of FSM)

* If BMM 0: record time

* If BMM 1 and changed or BMM 0 and changed: capture dout_0 = din_0, capture dout_1 = time delta


* Record Fifo occupancy changes

* byte mask/match 0 on din.data0[8;8] == 8b_00000000

* byte mask/match 1 on din.data0[8;8] == 8b_SSSSSSSS

* byte mask/match 2 on din.data0[8;16] == 8b_xx000000

* byte mask/match 3 on din.data0[8;16] == 8b_xxSSSSSS

* If BMM 0 changed or BMM 1 changed or BMM 2 changed or BMM 3 changed: capture dout_0 = din_0


* Two independent traces

* byte mask/match 0 on din.data0[8;0] == 8b_xxx00xxx

* byte mask/match 1 on din.data1[8;24] == 8b_xx11xxxx

* If BMM 0: capture dout_0 = d0_data,

* If BMM 1 and changed : capture dout_1 = d1_data


"""

{
    /*b Default clock and reset
     */
    default clock clk;
    default reset active_low reset_n;

    /*b State and combs */
    clocked t_timer_state timer_state = {*=0};
    clocked t_recorded_state recorded_state = {*=0};
    clocked t_analyzer_data4[5] data = {*=0};

    comb t_analyzer_data4 pretrigger_data;
    comb t_match_combs match_combs;
    net bit[8][4] match_conds;

    comb t_analyzer_trigger_cfg_data_source[2] trigger_cfg_ds;
    
    clocked bit[32][2] data_out = {*=0};
    clocked  t_analyzer_trace_op4 trace_op ={*=0};

    comb t_analyzer_trigger_cfg_data_action[2] trigger_cfg_m;

    /*b Timer value state
     */
    timer_value_logic "Timer value logic": {
        full_switch (trigger_cfg.timer_div) {
        case 2b00: {
            timer_state.value <= timer_value.value[32;0];
        }
        case 2b01: {
            timer_state.value <= timer_value.value[32;8];
        }
        case 2b10: {
            timer_state.value <= timer_value.value[32;16];
        }
        case 2b11: {
            timer_state.value <= timer_value.value[32;24];
        }
        }

        if (!trigger_cfg.enable) {
            timer_state <= timer_state;
        }
    }

    /*b Pretrigger data stage, record incoming data and implement 'only valid if changing'
     */
    pretrigger_data "Pretrigger data stage": {
        // data[0] is data in to byte mask match
        //
        // data[1] aligns with output of byte mask match, match_conds
        //
        // data[2] aligns with matched[] = output of analyzer_trigger_simple_byte
        //
        // data[3] aligns with dds_set_0/1

        if (din.valid || data[0].valid) {
            data[0].valid <= 0;
            if (trigger_cfg.enable) {
                data[0] <= din;
            }
        }

        if (data[0].valid || data[1].valid) {
            data[1].valid <= 0;
            if (data[0].valid) {
                data[1] <= data[0];
            }
        }

        pretrigger_data = data[0];

        if (data[1].valid || data[2].valid) {
            data[2].valid <= 0;
            if (data[1].valid) {
                data[2] <= data[1];
            }
        }

        if (data[2].valid || data[3].valid) {
            data[3].valid <= 0;
            if (data[2].valid) {
                data[3] <= data[2];
            }
        }

        match_combs.data = data[3];
        match_combs.data_changing = 0;

        if (data[3].data_0 != data[2].data_0) {
            match_combs.data_changing = 1;
        }
        if (data[3].data_1 != data[2].data_1) {
            match_combs.data_changing = 1;
        }
        if (data[3].data_2 != data[2].data_2) {
            match_combs.data_changing = 1;
        }
        if (data[3].data_3 != data[2].data_3) {
            match_combs.data_changing = 1;
        }

    }

    /*b Trigger byte matching and combining
     */
    trigger_byte "Trigger byte matching": {

        analyzer_trigger_simple_byte t0( clk <- clk, reset_n <= reset_n,
                                         din <= pretrigger_data,
                                         match_conds => match_conds[0],
                                         trigger_cfg_byte <= trigger_cfg.tb_0);
        analyzer_trigger_simple_byte t1( clk <- clk, reset_n <= reset_n,
                                         din <= pretrigger_data,
                                         match_conds => match_conds[1],
                                         trigger_cfg_byte <= trigger_cfg.tb_1);
        analyzer_trigger_simple_byte t2( clk <- clk, reset_n <= reset_n,
                                         din <= pretrigger_data,
                                         match_conds => match_conds[2],
                                         trigger_cfg_byte <= trigger_cfg.tb_2);
        analyzer_trigger_simple_byte t3( clk <- clk, reset_n <= reset_n,
                                         din <= pretrigger_data,
                                         match_conds => match_conds[3],
                                         trigger_cfg_byte <= trigger_cfg.tb_3);

        trigger_cfg_m[0] = trigger_cfg.data_action_0;
        trigger_cfg_m[1] = trigger_cfg.data_action_1;
        match_combs.matched = 0;
        if (match_combs.data.valid) {
            for (m; 2) {
                match_combs.matched[m] = (
                    match_conds[0][trigger_cfg_m[m].cond_0] &
                    match_conds[1][trigger_cfg_m[m].cond_1] &
                    match_conds[2][trigger_cfg_m[m].cond_2] &
                    match_conds[3][trigger_cfg_m[m].cond_3]
                    );
            }
        }

        match_combs.record_time = 0;
        match_combs.record_data = 0;
        match_combs.capture_data = 0;
        if (match_combs.matched[0] && (!trigger_cfg.data_action_0.only_if_changing || match_combs.data_changing)) {
            match_combs.record_time |= trigger_cfg.data_action_0.record_time;
            match_combs.record_data |= trigger_cfg.data_action_0.record_data;
            match_combs.capture_data |= trigger_cfg.data_action_0.capture_data;
        }
        if (match_combs.matched[1] && (!trigger_cfg.data_action_1.only_if_changing || match_combs.data_changing)) {
            match_combs.record_time |= trigger_cfg.data_action_1.record_time;
            match_combs.record_data |= trigger_cfg.data_action_1.record_data;
            match_combs.capture_data |= trigger_cfg.data_action_1.capture_data;
        }

    }

    /*b Data output generation (and recording for deltas)
     */
    data_out_generation "Data out generation": {
        trigger_cfg_ds[0] = trigger_cfg.data_source_0;
        trigger_cfg_ds[1] = trigger_cfg.data_source_1;
        trace_op.capture <= 0;
        for (i; 2) {
            if (match_combs.capture_data[i]) {
                trace_op.capture[i] <= 1;
                full_switch (trigger_cfg_ds[i]) {
                case atc_data_source_din_0: {
                    data_out[i] <= match_combs.data.data_0;
                }
                case atc_data_source_din_1: {
                    data_out[i] <= match_combs.data.data_1;
                }
                case atc_data_source_timer: {
                    data_out[i] <= timer_state.value;
                }
                case atc_data_source_timer_delta: {
                    data_out[i] <= timer_state.value - recorded_state.timer;
                }
                }
            }
        }
        if (match_combs.record_time) {
            recorded_state.timer <= timer_state.value;
        }
        if (match_combs.record_data) {
            recorded_state.data[0] <= match_combs.data.data_0;
            recorded_state.data[1] <= match_combs.data.data_1;
        }
        dout.valid = 0;
        dout.data_0 = data_out[0];
        dout.data_1 = data_out[1];
        dout.data_2 = 0; // data_out[2];
        dout.data_3 = 0; // data_out[3];
    }
    
    /*b Done
     */
}
